`timescale 1ps/1ps

#define SEED_SIZE 512 // 64*8

module ExpandS_tb;
    //Parameters match DUT
    localparam K = 8;
    localparam L = 7;
    localparam N = 256;
    localparam ETA = 2;                                 
    localparam COEFF_WIDTH = 4;          
    localparam DATA_IN_BITS = 64;        
    localparam DATA_OUT_BITS = 64;
    
    //DUT signals
    logic                             clk, rst, start, done;
    logic [`SEED_SIZE-1 : 0]          rho;
    logic [COEFF_WIDTH * N - 1 : 0]   s1[L];
    logic [COEFF_WIDTH * N - 1 : 0]   s2[K];

    // Instantiate the DUT
    ExpandS #(
        .K(K),
        .L(L),
        .N(N),
        .ETA(ETA),
        .COEFF_WIDTH(COEFF_WIDTH),
        .DATA_IN_BITS(DATA_IN_BITS),
        .DATA_OUT_BITS(DATA_OUT_BITS)
    ) dut (
        .clk(clk),
        .rst(rst),
        .start(start),
        .rho(rho),
        .done(done),
        .s1(s1),
        .s2(s2)
    );

    // Test instance
    initial clk = 0;
    always #5 clk = ~clk;

    initial begin
        rst = 1; 
        repeat (5) @(posedge clk);
        rst = 0;
    end

    initial begin
        //wait for reset to complete
        wait (!rst);
        repeat (5) @(posedge clk);

        //pulse start and push data in
        @(posedge clk);
        start = 1;
        // =================== WRITE YOUR TEST INPUT HERE ===================
        rho = 512'h
                1234567890abcdef_1234567890abcdef_
                1234567890abcdef_1234567890abcdef_
                1234567890abcdef_1234567890abcdef_
                1234567890abcdef_1234567890abcdef;
        @(posedge clk);
        start = 0;

        //wait for operation to complete
        wait(done);
        @(posedge clk);
        $write("s1 = ");
        foreach (s1[i]) $write("0x%0h ", s1[i]);
        $write("\n");
                  
        $write("s2 = ");
        foreach (s2[i]) $write("0x%0h ", s2[i]);
        $write("\n");
        #50 $finish;
    end
endmodule