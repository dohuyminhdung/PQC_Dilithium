`timescale 1ns / 1ps
// Algorithm 7: Sign a Signature (see FIPS 204 page 25, slide 35)
// Deterministic algorithm to generate a signature for a formatted message M_
// Input: private key sk, formatted message M_, random seed rnd
// Output: signature si

module Sign_internal #(
)(
);
endmodule